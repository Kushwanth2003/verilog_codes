module clk_buf(input mclk,output bufclk);
	buf(bufclk,mclk);
endmodule

